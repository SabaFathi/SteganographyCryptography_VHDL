library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

use work.AES_DEPENDENCY_PKG.ALL;

entity column_mixer is
port(in_matrix : in matrix_4X4;

	  clk : in std_logic;
	  enable : in std_logic;

	  out_matrix : out matrix_4X4);
end column_mixer;

architecture Behavioral of column_mixer is
begin

	process(clk)
	variable helper_vector : std_logic_vector(7 downto 0);
	variable helper_vector2 : std_logic_vector(7 downto 0);
	variable helper_vector3 : std_logic_vector(7 downto 0);
	variable helper_vector4 : std_logic_vector(7 downto 0);
	variable helper_carry1 : std_logic_vector(8 downto 0);
	variable helper_carry2 : std_logic_vector(8 downto 0);
	begin
		if(rising_edge(clk))
		then
			if(enable = '1')
			then
				--for each column:
				-- | 2 3 1 1 |          | c0 |   | 2*c0 + 3*c1 + 1*c2 + 1* c3 |
				-- | 1 2 3 1 | multiply | c1 | = | 1*c0 + 2*c1 + 3*c2 + 1* c3 |
				-- | 1 1 2 3 |          | c2 |   | 1*c0 + 1*c1 + 2*c2 + 3* c3 |
				-- | 3 1 1 2 |          | c3 |   | 3*c0 + 1*c1 + 1*c2 + 2* c3 |
				
				--GALOIS_FIELD_L_TABLE(02) = X"19"
				--GALOIS_FIELD_L_TABLE(03) = X"01"
				
				--column 0:
				helper_vector  := in_matrix(0, 0);
				helper_vector2 := in_matrix(1, 0);
				helper_vector3 := in_matrix(2, 0);
				helper_vector4 := in_matrix(3, 0);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"01";
				out_matrix(0, 0) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8)))) --add with carry
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector3)
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"01";
				out_matrix(1, 0) <= (helper_vector)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"01";
				out_matrix(2, 0) <= (helper_vector)
										 XOR (helper_vector2)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"01";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"19";
				out_matrix(3, 0) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (helper_vector2)
										 XOR (helper_vector3)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				--column 1:
				helper_vector  := in_matrix(0, 1);
				helper_vector2 := in_matrix(1, 1);
				helper_vector3 := in_matrix(2, 1);
				helper_vector4 := in_matrix(3, 1);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"01";
				out_matrix(0, 1) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector3)
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"01";
				out_matrix(1, 1) <= (helper_vector)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"01";
				out_matrix(2, 1) <= (helper_vector)
										 XOR (helper_vector2)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"01";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"19";
				out_matrix(3, 1) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (helper_vector2)
										 XOR (helper_vector3)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				--column 2:
				helper_vector  := in_matrix(0, 2);
				helper_vector2 := in_matrix(1, 2);
				helper_vector3 := in_matrix(2, 2);
				helper_vector4 := in_matrix(3, 2);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"01";
				out_matrix(0, 2) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector3)
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"01";
				out_matrix(1, 2) <= (helper_vector)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"01";
				out_matrix(2, 2) <= (helper_vector)
										 XOR (helper_vector2)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"01";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"19";
				out_matrix(3, 2) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (helper_vector2)
										 XOR (helper_vector3)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				--column 3:
				helper_vector  := in_matrix(0, 3);
				helper_vector2 := in_matrix(1, 3);
				helper_vector3 := in_matrix(2, 3);
				helper_vector4 := in_matrix(3, 3);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"01";
				out_matrix(0, 3) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector3)
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector2))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"01";
				out_matrix(1, 3) <= (helper_vector)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))))
										 XOR (helper_vector4);
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector3))) + X"19";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"01";
				out_matrix(2, 3) <= (helper_vector)
										 XOR (helper_vector2)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
				helper_carry1 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector))) + X"01";
				helper_carry2 := ('0' & GALOIS_FIELD_L_TABLE(conv_integer(helper_vector4))) + X"19";
				out_matrix(3, 3) <= (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry1(7 downto 0) + helper_carry1(8 downto 8))))
										 XOR (helper_vector2)
										 XOR (helper_vector3)
										 XOR (GALOIS_FIELD_E_TABLE(conv_integer(helper_carry2(7 downto 0) + helper_carry2(8 downto 8))));
				
			end if;
		end if;
	end process;

end Behavioral;
